`define module_name CORDIC_Top
`define ROTATE
`define PIPELINE
`define RADIAN_16
`define XY_BITS 17
`define THETA_BITS 17
`define ITERATIONS 16
`define ITERATION_BITS 4
